`define UTILS

module FF(clk, en, D, Q);
  parameter WIDTH = 1;
  parameter INIT  = 0;
 
  input wire                clk;
  input wire                en;
  input wire   [WIDTH-1:0]  D;
  output reg   [WIDTH-1:0]  Q = INIT;
  
  always @ (posedge clk) begin
    if(en) begin
      Q <= D;
    end
  end
endmodule
