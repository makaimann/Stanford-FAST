`define OPTIONS

// Data Integrity Scoreboard Options
//`define SB_SANITY
//`define EMBED
`define ARBITER

// FIFO Options
//`define SANITY
`define ARRAY

// DWRR Arbiter Options
`define COMB_UPDATE

// Parameters
`define FIFO_DEPTH 32
`define FIFO_DWIDTH 32
`define ARB_QWID 16
