`define OPTIONS

// Data Integrity Scoreboard Options
//`define SB_SANITY
//`define EMBED
//`define ARBITER

// FIFO Options
//`define SANITY
`define ARRAY

// DWRR Arbiter Options
//`define COMB_UPDATE

// Parameters
`define FIFO_DEPTH 8
`define FIFO_DWIDTH 8
`define ARB_QWID 8
