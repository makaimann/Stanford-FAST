`define OPTIONS

// Data Integrity Scoreboard Options
//`define SB_SANITY
//`define EMBED
`define ARBITER

// FIFO Options
//`define SANITY
//`define ARRAY

// DWRR Arbiter Options
`define COMB_UPDATE
